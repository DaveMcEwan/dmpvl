../usbFullSpeedSerial/driveHost.sv