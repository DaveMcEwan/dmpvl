.title PWM into Low-Pass Filter with optional LED
* Voltage source is o_pwm[i] driven by delta-sigma modulated 1.8V on GPIO.
* o_pwm pins may be low-pass filtered for sampling with oscilloscope.

* Unicode-schematics pallet: ─ │ ┌ ┐ ├ ┤ ┬ ┴ ┼ ⏚ Ω

.param jumperLpf=1 jumperLed=1

Vpin fpgaPin 0 dc 0 ac 1 PULSE (0 1.8 1u 10n 10n 0.208u 0.416u)
Vled ledCathode 0 dc 0 ; Ammeter
.if(jumperLpf && jumperLed)

  *   │           Vpin
  *   ├─fpgaPin───(+ 1.8V -)──────────────────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rlpf1                   Clpf1
  *   ├───[68Ω]───────lpfOut──────|100nF|─────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rprotect                  Dled                  Vled
  *   ├───[47Ω]───────ledAnode──────|>|─────ledCathode────(+ 0V -)────┐
  *   │                                                               ⏚

  Rlpf1 fpgaPin lpfOut 68
  Clpf1 lpfOut 0 100n
  Rprotect fpgaPin ledAnode 47
  Dled ledAnode ledCathode LED7030090

.elseif(jumperLed)

  *   │           Vpin
  *   ├─fpgaPin───(+ 1.8V -)──────────────────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rdummy                  Cdummy
  *   ├───[0Ω]────────lpfOut──────|0nF|───────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rprotect                  Dled                  Vled
  *   ├───[47Ω]───────ledAnode──────|>|─────ledCathode────(+ 0V -)────┐
  *   │                                                               ⏚

  Rdummy fpgaPin lpfOut 0
  Cdummy lpfOut 0 0
  Rprotect fpgaPin ledAnode 47
  Dled ledAnode ledCathode LED7030090

.elseif(jumperLpf)

  *   │           Vpin
  *   ├─fpgaPin───(+ 1.8V -)──────────────────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rlpf1                   Clpf1
  *   ├───[68Ω]───────lpfOut──────|100nF|─────────────────────────────┐
  *   │                                                               ⏚
  *   │
  *   │   Rdummy                    Cdummy                Vled
  *   ├───[0Ω]────────ledAnode──────|0nF|───ledCathode────(+ 0V -)────┐
  *   │                                                               ⏚

  Rlpf1 fpgaPin lpfOut 68
  Clpf1 lpfOut 0 100n
  Rdummy fpgaPin ledAnode 0
  Cdummy ledAnode ledCathode 0

.endif


* {{{ LED models

* Multicomp Pro 3mm Round LED Lamp, Red, AlGaAs/GaAs, 703-0090
* Vf=1.8V Vr=4V If=30mA trr=3uS
.MODEL LED7030090 D (
+ IS=93.2p RS=42m N=3.73
+ BV=4 IBV=10u
+ CJO=2.97P VJ=0.75 M=0.333
+ TT=4.32U)

*Typ RED GaAs LED: Vf=1.7V Vr=4V If=40mA trr=3uS
.MODEL LED1 D (IS=93.2P RS=42M N=3.73 BV=4 IBV=10U
+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)

*Typ RED,GREEN,YELLOW,AMBER GaAs LED: Vf=2.1V Vr=4V If=40mA trr=3uS
.MODEL LED2 D (IS=93.1P RS=42M N=4.61 BV=4 IBV=10U
+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)

*Typ BLUE SiC LED: Vf=3.4V Vr=5V If=40mA trr=3uS
.MODEL LED3 D (IS=93.1P RS=42M N=7.47 BV=5 IBV=30U
+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)

* }}} LED models


.control

** print
*set width=150
*set height=100k
*print col fpgaPin Vpin#branch lpfOut ledAnode Vled#branch > build/pwmFilter.foo.txt

** write
*set filetype=ascii
*write build/pwmFilter.foo.txt fpgaPin Vpin#branch lpfOut ledAnode Vled#branch

* wrdata
set wr_singlescale
set wr_vecnames

* plot,hardcopy
set hcopydevtype=postscript
set hcopypscolor = 0
set color0 = rgb:f/f/e ; Background
set color1 = rgb:0/0/0 ; Grid, Text
set color2 = rgb:0/0/0 ; fpgaPin, Voltage
set color3 = rgb:0/0/f ; Vpin#branch, Current
set color4 = rgb:0/f/0 ; lpfOut, Voltage
set color5 = rgb:f/0/0 ; ledAnode, Voltage
set color6 = rgb:8/8/8 ; Vled#branch, Current


tran 1n 30u
wrdata build/pwmFilter.tran.txt fpgaPin Vpin#branch lpfOut ledAnode Vled#branch
plot all
hardcopy build/pwmFilter.tran.ps fpgaPin Vpin#branch lpfOut ledAnode Vled#branch
+ ylimit -0.5 2.0


ac DEC 100 0.1kHz 1000kHz
wrdata build/pwmFilter.ac.txt fpgaPin Vpin#branch lpfOut ledAnode Vled#branch
plot all
hardcopy build/pwmFilter.ac.ps vdb(fpgaPin) vdb(Vpin#branch) vdb(lpfOut) vdb(ledAnode) vdb(Vled#branch)
set color2 = rgb:0/f/0 ; lpfOut, Voltage
hardcopy build/pwmFilter.ac.lpfOut.ps vdb(lpfOut)

quit
.endc

.end
