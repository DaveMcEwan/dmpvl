`include "dff.vh"

module corrCountLogdrop #(
  parameter DATA_W = 8,
  parameter TIME_W = 8
) (
  input wire                i_clk,
  input wire                i_rst,
  input wire                i_cg,

  input  wire               i_x,
  input  wire               i_y,

  output wire [DATA_W-1:0]  o_countX,
  output wire [DATA_W-1:0]  o_countY,
  output wire [DATA_W-1:0]  o_countIsect,   // x AND y
  output wire [DATA_W-1:0]  o_countSymdiff, // x XOR y

  input  wire               i_tUpdate, // 1->Beginning of new window.
  input  wire [TIME_W-1:0]  i_tValue, // Initial value for t in this window.
  output wire [TIME_W-1:0]  o_t
);

`dff_cg_srst(reg [TIME_W-1:0], t, i_clk, i_cg, i_rst)
always @* t_d = i_tUpdate ? i_tValue : t_q + 1;

wire [DATA_W-1:0] incrValue;
logdropWindow #(
  .DATA_W         (DATA_W),
  .WINLEN         (1 << TIME_W),
  .ABSTRACT_MODEL (0)
) u_win (
  .i_t  (t_q),
  .i_x  ({DATA_W{1'b1}}),
  .o_y  (incrValue)
);

`dff_cg_srst(reg [DATA_W-1:0], countX, i_clk, i_cg, i_rst || i_tUpdate)
always @* countX_d = i_x ? countX_q + incrValue : countX_q;

`dff_cg_srst(reg [DATA_W-1:0], countY, i_clk, i_cg, i_rst || i_tUpdate)
always @* countY_d = i_y ? countY_q + incrValue : countY_q;

`dff_cg_srst(reg [DATA_W-1:0], countIsect, i_clk, i_cg, i_rst || i_tUpdate)
always @* countIsect_d = (i_x & i_y) ? countIsect_q + incrValue : countIsect_q;

`dff_cg_srst(reg [DATA_W-1:0], countSymdiff, i_clk, i_cg, i_rst || i_tUpdate)
always @* countSymdiff_d = (i_x ^ i_y) ? countSymdiff_q + incrValue : countSymdiff_q;

assign o_countX       = countX_q;
assign o_countY       = countY_q;
assign o_countIsect   = countIsect_q;
assign o_countSymdiff = countSymdiff_q;

endmodule
