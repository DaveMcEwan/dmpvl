../correlator/correlator.sv