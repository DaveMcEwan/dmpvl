// Stub to infer PS7.
(* X_CORE_INFO = "processing_system7_v5_5_processing_system7,Vivado 2017.3" *)
module ps7_ip (
  TTC0_WAVE0_OUT,
  TTC0_WAVE1_OUT,
  TTC0_WAVE2_OUT,

  USB0_PORT_INDCTL,
  USB0_VBUS_PWRSELECT,
  USB0_VBUS_PWRFAULT,

  // {{{ AXI GP0
  M_AXI_GP0_ARVALID,
  M_AXI_GP0_AWVALID,
  M_AXI_GP0_BREADY,
  M_AXI_GP0_RREADY,
  M_AXI_GP0_WLAST,
  M_AXI_GP0_WVALID,
  M_AXI_GP0_ARID,
  M_AXI_GP0_AWID,
  M_AXI_GP0_WID,
  M_AXI_GP0_ARBURST,
  M_AXI_GP0_ARLOCK,
  M_AXI_GP0_ARSIZE,
  M_AXI_GP0_AWBURST,
  M_AXI_GP0_AWLOCK,
  M_AXI_GP0_AWSIZE,
  M_AXI_GP0_ARPROT,
  M_AXI_GP0_AWPROT,
  M_AXI_GP0_ARADDR,
  M_AXI_GP0_AWADDR,
  M_AXI_GP0_WDATA,
  M_AXI_GP0_ARCACHE,
  M_AXI_GP0_ARLEN,
  M_AXI_GP0_ARQOS,
  M_AXI_GP0_AWCACHE,
  M_AXI_GP0_AWLEN,
  M_AXI_GP0_AWQOS,
  M_AXI_GP0_WSTRB,
  M_AXI_GP0_ACLK,
  M_AXI_GP0_ARREADY,
  M_AXI_GP0_AWREADY,
  M_AXI_GP0_BVALID,
  M_AXI_GP0_RLAST,
  M_AXI_GP0_RVALID,
  M_AXI_GP0_WREADY,
  M_AXI_GP0_BID,
  M_AXI_GP0_RID,
  M_AXI_GP0_BRESP,
  M_AXI_GP0_RRESP,
  M_AXI_GP0_RDATA,
  // }}} AXI GP0

  // {{{ AXI GP1
  M_AXI_GP1_ARVALID,
  M_AXI_GP1_AWVALID,
  M_AXI_GP1_BREADY,
  M_AXI_GP1_RREADY,
  M_AXI_GP1_WLAST,
  M_AXI_GP1_WVALID,
  M_AXI_GP1_ARID,
  M_AXI_GP1_AWID,
  M_AXI_GP1_WID,
  M_AXI_GP1_ARBURST,
  M_AXI_GP1_ARLOCK,
  M_AXI_GP1_ARSIZE,
  M_AXI_GP1_AWBURST,
  M_AXI_GP1_AWLOCK,
  M_AXI_GP1_AWSIZE,
  M_AXI_GP1_ARPROT,
  M_AXI_GP1_AWPROT,
  M_AXI_GP1_ARADDR,
  M_AXI_GP1_AWADDR,
  M_AXI_GP1_WDATA,
  M_AXI_GP1_ARCACHE,
  M_AXI_GP1_ARLEN,
  M_AXI_GP1_ARQOS,
  M_AXI_GP1_AWCACHE,
  M_AXI_GP1_AWLEN,
  M_AXI_GP1_AWQOS,
  M_AXI_GP1_WSTRB,
  M_AXI_GP1_ACLK,
  M_AXI_GP1_ARREADY,
  M_AXI_GP1_AWREADY,
  M_AXI_GP1_BVALID,
  M_AXI_GP1_RLAST,
  M_AXI_GP1_RVALID,
  M_AXI_GP1_WREADY,
  M_AXI_GP1_BID,
  M_AXI_GP1_RID,
  M_AXI_GP1_BRESP,
  M_AXI_GP1_RRESP,
  M_AXI_GP1_RDATA,
  // }}} AXI GP1

  FCLK_CLK0,
  FCLK_RESET0_N,

  MIO,

  // {{{ DDR
  DDR_CAS_n,
  DDR_CKE,
  DDR_Clk_n,
  DDR_Clk,
  DDR_CS_n,
  DDR_DRSTB,
  DDR_ODT,
  DDR_RAS_n,
  DDR_WEB,
  DDR_BankAddr,
  DDR_Addr,
  DDR_VRN,
  DDR_VRP,
  DDR_DM,
  DDR_DQ,
  DDR_DQS_n,
  DDR_DQS,
  // }}} DDR

  PS_SRSTB,
  PS_CLK,
  PS_PORB
)

/* synthesis syn_black_box black_box_pad_pin="TTC0_WAVE0_OUT,TTC0_WAVE1_OUT,TTC0_WAVE2_OUT,USB0_PORT_INDCTL[1:0],USB0_VBUS_PWRSELECT,USB0_VBUS_PWRFAULT,M_AXI_GP0_ARVALID,M_AXI_GP0_AWVALID,M_AXI_GP0_BREADY,M_AXI_GP0_RREADY,M_AXI_GP0_WLAST,M_AXI_GP0_WVALID,M_AXI_GP0_ARID[11:0],M_AXI_GP0_AWID[11:0],M_AXI_GP0_WID[11:0],M_AXI_GP0_ARBURST[1:0],M_AXI_GP0_ARLOCK[1:0],M_AXI_GP0_ARSIZE[2:0],M_AXI_GP0_AWBURST[1:0],M_AXI_GP0_AWLOCK[1:0],M_AXI_GP0_AWSIZE[2:0],M_AXI_GP0_ARPROT[2:0],M_AXI_GP0_AWPROT[2:0],M_AXI_GP0_ARADDR[31:0],M_AXI_GP0_AWADDR[31:0],M_AXI_GP0_WDATA[31:0],M_AXI_GP0_ARCACHE[3:0],M_AXI_GP0_ARLEN[3:0],M_AXI_GP0_ARQOS[3:0],M_AXI_GP0_AWCACHE[3:0],M_AXI_GP0_AWLEN[3:0],M_AXI_GP0_AWQOS[3:0],M_AXI_GP0_WSTRB[3:0],M_AXI_GP0_ACLK,M_AXI_GP0_ARREADY,M_AXI_GP0_AWREADY,M_AXI_GP0_BVALID,M_AXI_GP0_RLAST,M_AXI_GP0_RVALID,M_AXI_GP0_WREADY,M_AXI_GP0_BID[11:0],M_AXI_GP0_RID[11:0],M_AXI_GP0_BRESP[1:0],M_AXI_GP0_RRESP[1:0],M_AXI_GP0_RDATA[31:0],M_AXI_GP1_ARVALID,M_AXI_GP1_AWVALID,M_AXI_GP1_BREADY,M_AXI_GP1_RREADY,M_AXI_GP1_WLAST,M_AXI_GP1_WVALID,M_AXI_GP1_ARID[11:0],M_AXI_GP1_AWID[11:0],M_AXI_GP1_WID[11:0],M_AXI_GP1_ARBURST[1:0],M_AXI_GP1_ARLOCK[1:0],M_AXI_GP1_ARSIZE[2:0],M_AXI_GP1_AWBURST[1:0],M_AXI_GP1_AWLOCK[1:0],M_AXI_GP1_AWSIZE[2:0],M_AXI_GP1_ARPROT[2:0],M_AXI_GP1_AWPROT[2:0],M_AXI_GP1_ARADDR[31:0],M_AXI_GP1_AWADDR[31:0],M_AXI_GP1_WDATA[31:0],M_AXI_GP1_ARCACHE[3:0],M_AXI_GP1_ARLEN[3:0],M_AXI_GP1_ARQOS[3:0],M_AXI_GP1_AWCACHE[3:0],M_AXI_GP1_AWLEN[3:0],M_AXI_GP1_AWQOS[3:0],M_AXI_GP1_WSTRB[3:0],M_AXI_GP1_ACLK,M_AXI_GP1_ARREADY,M_AXI_GP1_AWREADY,M_AXI_GP1_BVALID,M_AXI_GP1_RLAST,M_AXI_GP1_RVALID,M_AXI_GP1_WREADY,M_AXI_GP1_BID[11:0],M_AXI_GP1_RID[11:0],M_AXI_GP1_BRESP[1:0],M_AXI_GP1_RRESP[1:0],M_AXI_GP1_RDATA[31:0],FCLK_CLK0,FCLK_RESET0_N,MIO[53:0],DDR_CAS_n,DDR_CKE,DDR_Clk_n,DDR_Clk,DDR_CS_n,DDR_DRSTB,DDR_ODT,DDR_RAS_n,DDR_WEB,DDR_BankAddr[2:0],DDR_Addr[14:0],DDR_VRN,DDR_VRP,DDR_DM[3:0],DDR_DQ[31:0],DDR_DQS_n[3:0],DDR_DQS[3:0],PS_SRSTB,PS_CLK,PS_PORB" */;
  output        TTC0_WAVE0_OUT;
  output        TTC0_WAVE1_OUT;
  output        TTC0_WAVE2_OUT;

  output [1:0]  USB0_PORT_INDCTL;
  output        USB0_VBUS_PWRSELECT;
  input         USB0_VBUS_PWRFAULT;

  // {{{ GP0
  output        M_AXI_GP0_ARVALID;
  output        M_AXI_GP0_AWVALID;
  output        M_AXI_GP0_BREADY;
  output        M_AXI_GP0_RREADY;
  output        M_AXI_GP0_WLAST;
  output        M_AXI_GP0_WVALID;
  output [11:0] M_AXI_GP0_ARID;
  output [11:0] M_AXI_GP0_AWID;
  output [11:0] M_AXI_GP0_WID;
  output [1:0]  M_AXI_GP0_ARBURST;
  output [1:0]  M_AXI_GP0_ARLOCK;
  output [2:0]  M_AXI_GP0_ARSIZE;
  output [1:0]  M_AXI_GP0_AWBURST;
  output [1:0]  M_AXI_GP0_AWLOCK;
  output [2:0]  M_AXI_GP0_AWSIZE;
  output [2:0]  M_AXI_GP0_ARPROT;
  output [2:0]  M_AXI_GP0_AWPROT;
  output [31:0] M_AXI_GP0_ARADDR;
  output [31:0] M_AXI_GP0_AWADDR;
  output [31:0] M_AXI_GP0_WDATA;
  output [3:0]  M_AXI_GP0_ARCACHE;
  output [3:0]  M_AXI_GP0_ARLEN;
  output [3:0]  M_AXI_GP0_ARQOS;
  output [3:0]  M_AXI_GP0_AWCACHE;
  output [3:0]  M_AXI_GP0_AWLEN;
  output [3:0]  M_AXI_GP0_AWQOS;
  output [3:0]  M_AXI_GP0_WSTRB;
  input         M_AXI_GP0_ACLK;
  input         M_AXI_GP0_ARREADY;
  input         M_AXI_GP0_AWREADY;
  input         M_AXI_GP0_BVALID;
  input         M_AXI_GP0_RLAST;
  input         M_AXI_GP0_RVALID;
  input         M_AXI_GP0_WREADY;
  input  [11:0] M_AXI_GP0_BID;
  input  [11:0] M_AXI_GP0_RID;
  input  [1:0]  M_AXI_GP0_BRESP;
  input  [1:0]  M_AXI_GP0_RRESP;
  input  [31:0] M_AXI_GP0_RDATA;
  // }}} GP0

  // {{{ GP1
  output        M_AXI_GP1_ARVALID;
  output        M_AXI_GP1_AWVALID;
  output        M_AXI_GP1_BREADY;
  output        M_AXI_GP1_RREADY;
  output        M_AXI_GP1_WLAST;
  output        M_AXI_GP1_WVALID;
  output [11:0] M_AXI_GP1_ARID;
  output [11:0] M_AXI_GP1_AWID;
  output [11:0] M_AXI_GP1_WID;
  output [1:0]  M_AXI_GP1_ARBURST;
  output [1:0]  M_AXI_GP1_ARLOCK;
  output [2:0]  M_AXI_GP1_ARSIZE;
  output [1:0]  M_AXI_GP1_AWBURST;
  output [1:0]  M_AXI_GP1_AWLOCK;
  output [2:0]  M_AXI_GP1_AWSIZE;
  output [2:0]  M_AXI_GP1_ARPROT;
  output [2:0]  M_AXI_GP1_AWPROT;
  output [31:0] M_AXI_GP1_ARADDR;
  output [31:0] M_AXI_GP1_AWADDR;
  output [31:0] M_AXI_GP1_WDATA;
  output [3:0]  M_AXI_GP1_ARCACHE;
  output [3:0]  M_AXI_GP1_ARLEN;
  output [3:0]  M_AXI_GP1_ARQOS;
  output [3:0]  M_AXI_GP1_AWCACHE;
  output [3:0]  M_AXI_GP1_AWLEN;
  output [3:0]  M_AXI_GP1_AWQOS;
  output [3:0]  M_AXI_GP1_WSTRB;
  input         M_AXI_GP1_ACLK;
  input         M_AXI_GP1_ARREADY;
  input         M_AXI_GP1_AWREADY;
  input         M_AXI_GP1_BVALID;
  input         M_AXI_GP1_RLAST;
  input         M_AXI_GP1_RVALID;
  input         M_AXI_GP1_WREADY;
  input  [11:0] M_AXI_GP1_BID;
  input  [11:0] M_AXI_GP1_RID;
  input  [1:0]  M_AXI_GP1_BRESP;
  input  [1:0]  M_AXI_GP1_RRESP;
  input  [31:0] M_AXI_GP1_RDATA;
  // }}} GP1

  output        FCLK_CLK0;
  output        FCLK_RESET0_N;

  inout  [53:0] MIO;

  // {{{ DDR
  inout         DDR_CAS_n;
  inout         DDR_CKE;
  inout         DDR_Clk_n;
  inout         DDR_Clk;
  inout         DDR_CS_n;
  inout         DDR_DRSTB;
  inout         DDR_ODT;
  inout         DDR_RAS_n;
  inout         DDR_WEB;
  inout  [2:0]  DDR_BankAddr;
  inout  [14:0] DDR_Addr;
  inout         DDR_VRN;
  inout         DDR_VRP;
  inout  [3:0]  DDR_DM;
  inout  [31:0] DDR_DQ;
  inout  [3:0]  DDR_DQS_n;
  inout  [3:0]  DDR_DQS;
  // }}} DDR

  inout         PS_SRSTB;
  inout         PS_CLK;
  inout         PS_PORB;
endmodule
