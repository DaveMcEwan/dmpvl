// USB spec r1.0

// Transition states.
// {d+, d-}
localparam LINE_SE0  = 2'b00; // Single-ended 0
localparam LINE_SE1  = 2'b11; // Single-ended 1
localparam LINE_J   = 2'b10; // Differential J
localparam LINE_K   = 2'b01; // Differential K


/*
7.1.6 Bit Stuffing
In order to ensure adequate signal transitions, bit stuffing is employed by the
transmitting device when sending a packet on the USB (see Figure 7-13 and
Figure 7-14).
A 0 is inserted after every six consecutive 1’s in the data stream before the
data is NRZI encoded to force a transition in the NRZI data stream.
This gives the receiver logic a data transition at least once every seven bit
times to guarantee the data and clock lock.
The receiver must decode the NRZI data, recognize the stuffed bits, and discard
them.
Bit stuffing is enabled beginning with the Sync Pattern and throughout the
entire transmission.
The data “one” that ends the Sync Pattern is counted as the first one in a
sequence.
Bit stuffing is always enforced, without exception.
If required by the bit stuffing rules, a zero bit will be inserted even if it
is the last bit before the end-of-packet (EOP) signal.
*/
localparam NRZI_MAXRL_ONES = 6;
localparam NRZI_ENC0_A = {LINE_J, LINE_K};
localparam NRZI_ENC0_B = {LINE_K, LINE_J};
localparam NRZI_ENC1_A = {LINE_K, LINE_K};
localparam NRZI_ENC1_B = {LINE_J, LINE_J};


/*
7.1.7 Sync Pattern
The NRZI bit pattern shown in Figure 7-15 is used as a synchronization pattern
and is prefixed to each
packet.
This pattern is equivalent to a data pattern of seven 0s followed by a 1.

8.2 SYNC Field, p145
All packets begin with a synchronization (SYNC) field, which is a coded
sequence that generates a maximum edge transition density.
The SYNC field appears on the bus as IDLE followed by the binary string
“KJKJKJKK”, in its NRZI encoding.
It is used by the input circuitry to align incoming data with the local clock
and is defined to be eight bits in length.
SYNC serves only as a synchronization mechanism and is not shown in the
following packet diagrams (refer to Section 7.1.7).
The last two bits in the SYNC field are a marker that is used to identify the
first bit of the PID.
All subsequent bits in the packet must be indexed from this point.
*/
// NOTE: A receiver can pinpoint SOP/PID by detecting only the last 3
// transitions (JKK)
// NOTE: Arranged LSB first, like all other data.
localparam SYNC_SOP = 8'b10000000;


/*
8.3.1 Packet Identifier Field, p145
A packet identifier (PID) immediately follows the SYNC field of every USB
packet.
A PID consists of a four bit packet type field followed by a four-bit check
field as shown in Figure 8-1.
The PID indicates the type of packet and, by inference, the format of the
packet and the type of error detection applied to the packet.
The four-bit check field of the PID insures reliable decoding of the PID so
that the remainder of the packet is interpreted correctly.
The PID check field is generated by performing a ones complement of the
packet type field.

The host and all functions must perform a complete decoding of all received PID
fields.
Any PID received with a failed check field or which decodes to a non-defined
value is assumed to be corrupted and it, as well as the remainder of the
packet, is ignored by the packet receiver.
If a function receives an otherwise valid PID for a transaction type or
direction that it does not support, the function must not respond.
For example, an IN only endpoint must ignore an OUT token.
PID types, codings, and descriptions are listed in Table 8-1.

PIDs are divided into four coding groups: TOKEN, DATA, HANDSHAKE, and SPECIAL,
with the first two transmitted PID bits (PID<1:0>) indicating which group.
This accounts for the distribution of PID codes.
*/
// {{{ Table 8-1 PID Types

// 2 LSBs determine coding group.
localparam PIDGROUP_TOKEN     = 2'b01;
localparam PIDGROUP_DATA      = 2'b11;
localparam PIDGROUP_HANDSHAKE = 2'b10;
localparam PIDGROUP_SPECIAL   = 2'b00;

// Address + endpoint number in host -> function transaction.
localparam PID_TOKEN_OUT = 4'b0001;

// Address + endpoint number in function -> host transaction.
localparam PID_TOKEN_IN = 4'b1001;

// Start of frame marker and frame number.
localparam PID_TOKEN_SOF = 4'b0101;

// Address + endpoint number in host -> function transaction for setup to a
// control endpoint.
localparam PID_TOKEN_SETUP = 4'b1101;

// Data packet PID even.
localparam PID_DATA_DATA0 = 4'b0011;

// Data packet PID odd.
localparam PID_DATA_DATA1 = 4'b1011;

// Data packet PID high-speed, high bandwidth isochronous transaction in a
// microframe (125us).
localparam PID_DATA_DATA2 = 4'b0111;

// Data packet PID high-speed for split and high bandwidth isochronous
// transactions
localparam PID_DATA_MDATA = 4'b1111;

// Receiver accepts error free data packet.
localparam PID_HANDSHAKE_ACK = 4'b0010;

// Receiving device cannot accept data or transmitting device cannot send data.
localparam PID_HANDSHAKE_NAK = 4'b1010;

// Endpoint is halted or a control pipe request is not supported.
localparam PID_HANDSHAKE_STALL = 4'b1110;

// No response yet from receiver.
localparam PID_HANDSHAKE_NYET = 4'b0110;

// (token) Host-issued preamble.
// Enables downstream bus traffic to low speed devices.
localparam PID_SPECIAL_PRE = 4'b1100;

// (handshake) Split Transaction Error Handshake (reuses PRE value).
localparam PID_SPECIAL_ERR = 4'b1100;

// (token) High-speed Split Transaction Token.
localparam PID_SPECIAL_SPLIT = 4'b1100;

// (token) High-speed flow control probe for a bulk/control endpoint.
localparam PID_SPECIAL_PING = 4'b0100;

// }}} Table 8-1 PID Types

/*
8.3.5.1 Token CRCs
A five-bit CRC field is provided for tokens and covers the ADDR and ENDP fields
of IN, SETUP, and OUT tokens or the time stamp field of an SOF token.
The generator polynomial is:
  G(x) = x^5 + x^2 + 1
The binary bit pattern that represents this polynomial is 00101.
If all token bits are received without error, the five-bit residual at the
receiver will be 01100 (x^4 + x^3).
*/
localparam TOKEN_CRC_POLYNOMIAL = 5'b00101;
localparam TOKEN_CRC_RESIDUAL = 5'b01100;

/*
8.3.5.2 Data CRCs
The data CRC is a 16-bit polynomial applied over the data field of a data
a packet.
The generating polynomial is:
  G(x) = x^16 + x^15 + x^2 + 1
The binary bit pattern that represents this polynomial is 1000000000000101.
If all data and CRC bits are received without error, the 16-bit residual will
be 1000000000001101.
*/
localparam DATA_CRC_POLYNOMIAL = 16'b1000000000000101;
localparam DATA_CRC_RESIDUAL = 16'b1000000000001101;

// 8.4.1 Token Packets          {PID:8b, ADDR:7b, ENDP:4b, CRC5:5b}
// 8.4.2 Start of Frame Packets {PID:8b, Frame Number:11b, CRC5:5b}
// 8.4.2 Data Packets           {PID:8b, data:0..1023b, CRC16:16b}
// 8.4.4 Handshake Packets      {PID:8b}
localparam TOKEN_FIELD_ADDR_LENGTH = 4'd7;
localparam TOKEN_FIELD_ENDP_LENGTH = 4'd4;
localparam SOF_FIELD_FRAMENUMBER_LENGTH = 4'd11;

// {{{ Table 9-4 Standard Request Codes

localparam BREQUEST_GET_STATUS        = 8'd0;
localparam BREQUEST_CLEAR_FEATURE     = 8'd1;
//localparam BREQUEST_reserved        = 8'd2;
localparam BREQUEST_SET_STATUS        = 8'd3;
//localparam BREQUEST_reserved        = 8'd4;
localparam BREQUEST_SET_ADDRESS       = 8'd5;
localparam BREQUEST_GET_DESCRIPTOR    = 8'd6;
localparam BREQUEST_SET_DESCRIPTOR    = 8'd7;
localparam BREQUEST_GET_CONFIGURATION = 8'd8;
localparam BREQUEST_SET_CONFIGURATION = 8'd9;
localparam BREQUEST_GET_INTERFACE     = 8'd10;
localparam BREQUEST_SET_INTERFACE     = 8'd11;
localparam BREQUEST_SYNCH_FRAME       = 8'd12;

localparam BREQUEST_CDC_SET = 8'h21;
localparam BREQUEST_CDC_GET = 8'h51;

// }}} Table 9-4 Standard Request Codes

// {{{ Table 9-5 Descriptor Types

localparam BDESCRIPTORTYPE_DEVICE         = 8'd1;
localparam BDESCRIPTORTYPE_CONFIGURATION  = 8'd2;
localparam BDESCRIPTORTYPE_STRING         = 8'd3;
localparam BDESCRIPTORTYPE_INTERFACE      = 8'd4;
localparam BDESCRIPTORTYPE_ENDPOINT       = 8'd5;
localparam BDESCRIPTORTYPE_DEVICEQUALIFIER = 8'd6;
localparam BDESCRIPTORTYPE_OTHERSPEED     = 8'd7;
localparam BDESCRIPTORTYPE_IFACEPOWER     = 8'd8;

localparam BDESCRIPTORTYPE_CS_INTERFACE   = 8'h24;

// }}} Table 9-5 Descriptor Types


// {{{ Defined Class Codes
// https://www.usb.org/defined-class-codes

localparam BASECLASS_UNKNOWN          = 8'h00; // Use class information in the Interface Descriptors
localparam BASECLASS_AUDIO            = 8'h01; // Audio
localparam BASECLASS_CDCCTRL          = 8'h02; // Communications and CDC Control
localparam BASECLASS_HID              = 8'h03; // Human Interface Device
localparam BASECLASS_PHYSICAL         = 8'h05; // Physical
localparam BASECLASS_IMAGE            = 8'h06; // Image
localparam BASECLASS_PRINTER          = 8'h07; // Printer
localparam BASECLASS_MASSSTORAGE      = 8'h08; // Mass Storage
localparam BASECLASS_HUB              = 8'h09; // Hub
localparam BASECLASS_CDCDATA          = 8'h0a; // CDC-Data
localparam BASECLASS_SMARTCARD        = 8'h0b; // Smart Card
localparam BASECLASS_CONTENTSECURITY  = 8'h0d; // Content Security
localparam BASECLASS_VIDEO            = 8'h0e; // Video
localparam BASECLASS_HEALTHCARE       = 8'h0f; // Personal Healthcare
localparam BASECLASS_AUDIOVIDEO       = 8'h10; // Audio/Video Devices
localparam BASECLASS_BILLBOARD        = 8'h11; // Billboard Device Class
localparam BASECLASS_CBRIDGE          = 8'h12; // USB Type-C Bridge Class
localparam BASECLASS_DIAGNOSTIC       = 8'hdc; // Diagnostic Device
localparam BASECLASS_WIRELESSCTRL     = 8'he0; // Wireless Controller
localparam BASECLASS_MISC             = 8'hef; // Miscellaneous
localparam BASECLASS_APPLICATION      = 8'hfe; // Application Specific
localparam BASECLASS_VENDOR           = 8'hff; // Vendor Specific

// }}} Defined Class Codes

localparam CDC_IFACE_SUBCLASS_DLCM  = 8'h01; // Direct Line Control Model
localparam CDC_IFACE_SUBCLASS_ACM   = 8'h02; // Abstract Control Model
localparam CDC_IFACE_SUBCLASS_TCM   = 8'h03; // Telephone Control Model
localparam CDC_IFACE_SUBCLASS_MCCM  = 8'h04; // Multi-Channel Control Model
localparam CDC_IFACE_SUBCLASS_CCM   = 8'h05; // CAPI Control Model
localparam CDC_IFACE_SUBCLASS_ENCM  = 8'h06; // Ethernet Networking Control Model
localparam CDC_IFACE_SUBCLASS_ANCM  = 8'h07; // ATM Networking Control Model

localparam ENDPTYPE_BULK       = 8'h02; // Bulk
localparam ENDPTYPE_INTERRUPT  = 8'h03; // Interrupt

// {{{ Table 13 bDescriptor SubType in Communications Class Functional Descriptors

// Header Functional Descriptor, which marks the beginning of the concatenated
// set of functional descriptors for the interface.
localparam BDESCRIPTORSUBTYPE_CDC_HEADER    = 8'h00;

// Call Management Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_CALLMGMT  = 8'h01;

// Abstract Control Management Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_ACM       = 8'h02;

// Direct Line Control Management Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_DLM       = 8'h03;

// Telephone Ringer Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_TR        = 8'h04;

// Telephone Call and Line State Reporting Capabilities Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_TC        = 8'h05;

// Union Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_UNION     = 8'h06;

// Country Selection Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_COUNTRY   = 8'h07;

// Telephone Operational Modes Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_TOM       = 8'h08;

// USB Terminal Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_USBTERM   = 8'h09;

// Network Channel Terminal Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_NETTERM   = 8'h0A;

// Protocol Unit Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_PU        = 8'h0B;

// Extension Unit Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_EU        = 8'h0C;

// Multi-Channel Management Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_MCM       = 8'h0D;

// CAPI Control Management Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_CAPICM    = 8'h0E;

// Ethernet Networking Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_ENET      = 8'h0F;

// ATM Networking Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_ATMNET    = 8'h10;

// Wireless Handset Control Model Functional Descriptor.
localparam BDESCRIPTORSUBTYPE_CDC_WHCM      = 8'h11;

// }}} Table 13 bDescriptor SubType in Communications Class Functional Descriptors
