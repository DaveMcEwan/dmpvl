../correlator/bpReg.sv