module example ();
  typedef struct packed {
    bit a;
    logic b;
    bit c;
  } foo;
endmodule
