../correlator/usbfsBpCorrelator.sv