`include "dff.vh"

module correlator #(
  parameter PRECISION = 20,
  parameter MAX_SAMPLE_RATE_NEGEXP = 15,
  parameter MAX_SAMPLE_JITTER_NEGEXP = 14
) (
  input wire          i_clk,
  input wire          i_rst,
  input wire          i_cg,

  input  wire         i_x,
  input  wire         i_y,

  input  wire [7:0]   i_bp_data,
  input  wire         i_bp_valid,
  output wire         o_bp_ready,

  output wire [7:0]   o_bp_data,
  output wire         o_bp_valid,
  input  wire         i_bp_ready
);

// maxWinLenExp is same as precision for accurate LogDrop window calculation.
localparam MAX_WINDOW_LENGTH_EXP = PRECISION;

genvar i;

wire [7:0]        pktfifo_o_data;
wire              pktfifo_o_empty;
wire              pktfifo_i_pop;

wire [$clog2(PRECISION)-1:0]                 windowLengthExp;
wire                                         windowShape;
wire [$clog2(MAX_SAMPLE_RATE_NEGEXP)-1:0]    sampleRateNegExp;
wire                                         sampleMode;
wire [$clog2(MAX_SAMPLE_JITTER_NEGEXP)-1:0]  sampleJitterNegExp;

bpReg #(
  .PRECISION                (PRECISION),
  .MAX_SAMPLE_RATE_NEGEXP   (MAX_SAMPLE_RATE_NEGEXP),
  .MAX_SAMPLE_JITTER_NEGEXP (MAX_SAMPLE_JITTER_NEGEXP)
) u_bpReg (
  .i_clk              (i_clk),
  .i_rst              (i_rst),
  .i_cg               (1'b1),

  .i_pktfifo_data   (pktfifo_o_data),
  .i_pktfifo_empty  (pktfifo_o_empty),
  .o_pktfifo_pop    (pktfifo_i_pop),

  .o_reg_windowLengthExp    (windowLengthExp),
  .o_reg_windowShape        (windowShape),
  .o_reg_sampleRateNegExp   (sampleRateNegExp),
  .o_reg_sampleMode         (sampleMode),
  .o_reg_sampleJitterNegExp (sampleJitterNegExp),

  .i_bp_data   (i_bp_data),
  .i_bp_valid  (i_bp_valid),
  .o_bp_ready  (o_bp_ready),

  .o_bp_data   (o_bp_data),
  .o_bp_valid  (o_bp_valid),
  .i_bp_ready  (i_bp_ready)
);

reg [7:0] pktfifo_i_data;
wire pktfifo_i_push = newWin || (pktIdx_q != 3'd0);
wire              _unused_pktfifo_o_full;
wire              _unused_pktfifo_o_pushed;
wire              _unused_pktfifo_o_popped;
wire [5:0]        _unused_pktfifo_o_wrptr;
wire [5:0]        _unused_pktfifo_o_rdptr;
wire [49:0]       _unused_pktfifo_o_valid;
wire [5:0]        _unused_pktfifo_o_nEntries;
wire [8*50-1:0]   _unused_pktfifo_o_entries;
fifo #(
  .WIDTH          (8),
  .DEPTH          (50),
  .FLOPS_NOT_MEM  (0)
) u_fifo (
  .i_clk      (i_clk),
  .i_rst      (i_rst),
  .i_cg       (1'b1),

  .i_flush    (1'b0), // TODO: Flush register for recovery.
  .i_push     (pktfifo_i_push),
  .i_pop      (pktfifo_i_pop),

  .i_data     (pktfifo_i_data),
  .o_data     (pktfifo_o_data),

  .o_empty    (pktfifo_o_empty),
  .o_full     (_unused_pktfifo_o_full),

  .o_pushed   (_unused_pktfifo_o_pushed),
  .o_popped   (_unused_pktfifo_o_popped),

  .o_wrptr    (_unused_pktfifo_o_wrptr),
  .o_rdptr    (_unused_pktfifo_o_rdptr),

  .o_valid    (_unused_pktfifo_o_valid),
  .o_nEntries (_unused_pktfifo_o_nEntries),

  .o_entries  (_unused_pktfifo_o_entries)
);

`dff_cg_srst(reg [MAX_WINDOW_LENGTH_EXP-1:0], t, i_clk, i_cg, i_rst, '0)
always @* t_d = newWin ? '0 : t_q + 1;

wire [MAX_WINDOW_LENGTH_EXP-1:0] tDoWrapVec;
generate for (i = 0; i < MAX_WINDOW_LENGTH_EXP; i=i+1) begin
  if (i == 0)
    assign tDoWrapVec[0] = (windowLengthExp == 0);
  else
    assign tDoWrapVec[i] = (windowLengthExp == i) && (&t_q[0 +: i]);
end endgenerate
wire newWin = |tDoWrapVec;

wire [MAX_WINDOW_LENGTH_EXP-1:0] rect_countX;
wire [MAX_WINDOW_LENGTH_EXP-1:0] rect_countY;
wire [MAX_WINDOW_LENGTH_EXP-1:0] rect_countIsect;
wire [MAX_WINDOW_LENGTH_EXP-1:0] rect_countSymdiff;
corrCountRect #(
  .TIME_W  (MAX_WINDOW_LENGTH_EXP)
) u_winRect (
  .i_clk          (i_clk),
  .i_rst          (i_rst),
  .i_cg           (1'b1),

  .i_x            (i_x),
  .i_y            (i_y),

  .o_countX       (rect_countX),
  .o_countY       (rect_countY),
  .o_countIsect   (rect_countIsect),
  .o_countSymdiff (rect_countSymdiff),

  .i_zeroCounts   (newWin)
);

// NOTE: Window coefficient is 1 sample out of of phase in order to meet timing.
// Therefore the X and Y inputs are also flopped.
// As winNum is pushed into the fifo before any results this is okay.
`dff_cg_norst(reg, x, i_clk, i_cg)
`dff_cg_norst(reg, y, i_clk, i_cg)
always @* y_d = i_y;
always @* x_d = i_x;

wire [PRECISION+MAX_WINDOW_LENGTH_EXP-1:0] logdrop_countX;
wire [PRECISION+MAX_WINDOW_LENGTH_EXP-1:0] logdrop_countY;
wire [PRECISION+MAX_WINDOW_LENGTH_EXP-1:0] logdrop_countIsect;
wire [PRECISION+MAX_WINDOW_LENGTH_EXP-1:0] logdrop_countSymdiff;
corrCountLogdrop #(
  .DATA_W  (PRECISION+MAX_WINDOW_LENGTH_EXP),
  .TIME_W  (MAX_WINDOW_LENGTH_EXP)
) u_winLogdrop (
  .i_clk          (i_clk),
  .i_rst          (i_rst),
  .i_cg           (1'b1),

  .i_x            (x_q),
  .i_y            (y_q),

  .o_countX       (logdrop_countX),
  .o_countY       (logdrop_countY),
  .o_countIsect   (logdrop_countIsect),
  .o_countSymdiff (logdrop_countSymdiff),

  .i_t            (t_q),
  .i_zeroCounts   (newWin)
);

// Wrapping window counter to be used only to check that packets have not been
// dropped.
`dff_upcounter(reg [7:0], winNum, i_clk, newWin, i_rst)

// Only the 8 most significant bits of the counters is reported
wire [7:0] pkt_countX = windowShape ?
  logdrop_countX[PRECISION+MAX_WINDOW_LENGTH_EXP-8 +: 8] :
  rect_countX[MAX_WINDOW_LENGTH_EXP-8 +: 8];

wire [7:0] pkt_countY = windowShape ?
  logdrop_countY[PRECISION+MAX_WINDOW_LENGTH_EXP-8 +: 8] :
  rect_countY[MAX_WINDOW_LENGTH_EXP-8 +: 8];

wire [7:0] pkt_countIsect = windowShape ?
  logdrop_countIsect[PRECISION+MAX_WINDOW_LENGTH_EXP-8 +: 8] :
  rect_countIsect[MAX_WINDOW_LENGTH_EXP-8 +: 8];

wire [7:0] pkt_countSymdiff = windowShape ?
  logdrop_countSymdiff[PRECISION+MAX_WINDOW_LENGTH_EXP-8 +: 8] :
  rect_countSymdiff[MAX_WINDOW_LENGTH_EXP-8 +: 8];

`dff_upcounter(reg [2:0], pktIdx, i_clk, pktfifo_i_push, i_rst || (pktIdx_q == 3'd4))

always @*
  case (pktIdx_q)
    3'd1:     pktfifo_i_data = pkt_countX;
    3'd2:     pktfifo_i_data = pkt_countY;
    3'd3:     pktfifo_i_data = pkt_countIsect;
    3'd4:     pktfifo_i_data = pkt_countSymdiff;
    default:  pktfifo_i_data = winNum_q;
  endcase

endmodule
