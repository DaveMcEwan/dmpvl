`ifndef AMBASPEC_SVH_
`define AMBASPEC_SVH_

localparam AXI_RESP_OKAY = 2'b00;
localparam AXI_RESP_EXOKAY = 2'b01; // Not supported in axi4lite
localparam AXI_RESP_SLVERR = 2'b10;
localparam AXI_RESP_DECERR = 2'b11;

`endif // AMBASPEC_SVH_
