../correlator/bpCorrelator.sv