module BUFG (
  input  wire         I,
  output wire         O
);

buf u0 (O, I);

endmodule
