module M;
  woops @(posedge clk) z = z - 1;
endmodule
